module memory();
integer memory[1023:0];
integer cache [3:0][7:0];
integer i;
    initial
    begin
        for (i=0; i<100; i=i+1)
        begin

        end

    end
endmodule